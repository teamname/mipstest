module driver();
  
  parameter D_ME = ""; //data mem
  parameter I_ME = ""; //instr mem
  parameter TEST_FILE = "";
  parameter TEST_SZ = 5;
  reg [9:0] inst_in;
  reg [7:0] data_in;
  reg [31:0] inst_out, data_out;
  reg clk, rst;
  
  integer k; //loop
  //test addr array
  reg [7:0] ins [TEST_SZ - 1:0];
  
  //expected output array
  reg [31:0] outs [TEST_SZ - 1:0]; 


  //file stuff
  integer file_handle,error,indx,num_bytes_in_line;
  reg [0:255] line_buffer;
  reg [639:0] err_str;
  
  forever #10 clk = ~clk; //create clock
  
  
  toplevel #(D_ME, I_ME) DUT (clk, rst, inst_in, data_in, inst_out, data_out); //instantiate module
  
  initial begin
    //initials
    clk = 1'b0;
    rst = 1'b1;
    data_in = 8'h00;
    inst_in = 10'h000;
    //setup test data from file
  file_handle = $fopen(TEST_FILE,?r?);
  error = $ferror(file_handle,err_str);
  if (error==0) begin
    for(k = 0; k < TEST_SZ*2 ; k = k+1)
      num_bytes_in_line = $fgets(line_buffer,file_handle);
      ins[k] = line_buffer;
      num_bytes_in_line = $fgets(line_buffer,file_handle);
      outs[k] = line_buffer;
    end 
  end
  else begin 
   $display(?Could not open file");
   $stop; 
  end

    #15 rst = 1'b0;
    #100000;
    
    for(k = 0; k < TEST_SZ; k = k + 1)
      data_in = ins[k];
      if(data_out != outs[k])
        $display("Unexpected output for k = %d, expected: %h, got : %h", k, outs[k], data_out);
      else
        $display("Output for k = %d was okay!", k); 
    end
    
    $stop;
  end //end initial
  
endmodule
