library verilog;
use verilog.vl_types.all;
entity exe is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        dummyE          : in     vl_logic;
        spriteE         : in     vl_logic;
        fontE           : in     vl_logic;
        backgroundE     : in     vl_logic;
        posE            : in     vl_logic;
        attrE           : in     vl_logic;
        visiE           : in     vl_logic;
        rd_E            : in     vl_logic_vector(4 downto 0);
        luiE            : in     vl_logic;
        md_start_E      : in     vl_logic;
        alu_out_sel     : in     vl_logic_vector(1 downto 0);
        forward_a_E     : in     vl_logic_vector(1 downto 0);
        forward_b_E     : in     vl_logic_vector(1 downto 0);
        alu_cnt_E       : in     vl_logic_vector(2 downto 0);
        src_a_E         : in     vl_logic_vector(31 downto 0);
        src_b_E         : in     vl_logic_vector(31 downto 0);
        data_in         : in     vl_logic_vector(31 downto 0);
        alu_out_M       : in     vl_logic_vector(31 downto 0);
        sign_imm_E      : in     vl_logic_vector(31 downto 0);
        pc_E            : in     vl_logic_vector(31 downto 0);
        src_b_out_E     : out    vl_logic_vector(31 downto 0);
        alu_out_E       : out    vl_logic_vector(31 downto 0);
        of_E            : out    vl_logic;
        md_run_E        : out    vl_logic;
        sprite_x        : out    vl_logic_vector(9 downto 0);
        sprite_y        : out    vl_logic_vector(8 downto 0);
        sprite_sel      : out    vl_logic_vector(4 downto 0);
        sprite_attr     : out    vl_logic;
        sprite_pos      : out    vl_logic;
        sprite_vis      : out    vl_logic;
        font_addr       : out    vl_logic_vector(10 downto 0);
        font_data       : out    vl_logic_vector(3 downto 0);
        font_en         : out    vl_logic;
        bck             : out    vl_logic_vector(1 downto 0);
        bck_ch_active   : out    vl_logic;
        font_ch_active  : out    vl_logic;
        font_clr        : out    vl_logic
    );
end exe;
